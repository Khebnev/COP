library IEEE;
use IEEE.std_logic_1164.all;

entity RGB_LED is
       port (
            
            );
end RGB_LED;
architecture communication of RGB_LED is
begin
        
end communication;