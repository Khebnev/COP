library IEEE;
use IEEE.std_logic_1164.all;

entity ControlBlock is
       port (  clk_enab: out std_logic; 
					clk: out std_logic;
					reset: out std_logic
            );
end ControlBlock;
architecture Ctrl of ControlBlock is
begin
        
end Ctrl;